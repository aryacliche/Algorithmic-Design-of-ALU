library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use Work; -- I forgot how to import the entity from another file

entity datapath is
	generic (
		INPUT_WIDTH: integer := 8;
		COUNTER_WIDTH: integer := 4
	);
	port (
		clk, t0, t1: in std_logic;
		p0: out std_logic; 
		a,b: in std_logic_vector (INPUT_WIDTH - 1 downto 0);
		p:   out std_logic_vector(2 * INPUT_WIDTH - 1 downto 0)
		);
end entity datapath;

architecture standard of datapath is
	
	-- component Add2 is  -- Adding the necessary components
	--    port (
	-- 		start: in std_logic; 
	-- 		done: out std_logic;
	-- 		A,B: in std_logic_vector (7 downto 0);
	-- 		C:   out std_logic_vector(7 downto 0);
	-- 		clk: in std_logic;
	-- 		reset: in std_logic);
	-- end component;

	signal ta : std_logic_vector(INPUT_WIDTH - 1 downto 0);
	signal t : std_logic_vector(INPUT_WIDTH * 2 downto 0);
	signal counter : unsigned(COUNTER_WIDTH - 1 downto 0);	-- Since we are only going to be using simple addition on it
	
	begin
		-- Structural stuff
		-- main_adder : Add2 port map(start, done, s1, s2, s3, clk, reset); 		-- Why is this adder so weird.
		
		p <= t(2 * INPUT_WIDTH - 1 downto 0); -- The output is connected to the t register (but we skip the MSB for some reason)
		p0 <= (AND (std_logic_vector(counter) xnor std_logic_vector(to_unsigned(INPUT_WIDTH, COUNTER_WIDTH)))); -- The predicate is the counter xor 8	(Has to be combinational logic therefore is outside of the process)

		process(clk, t0, t1)
		begin
			if rising_edge(clk) then
				if(t0 = '1') then -- We are in the reset state
					ta <= a;
					t <= (others => '0');
					counter <= (others => '0');
				
				elsif (t1 = '1') then -- We are in the LOOP_STATE part OR we just transitioned to DONE_STATE
					if(ta(0) = '1') then
						t(2 * INPUT_WIDTH downto INPUT_WIDTH) <= std_logic_vector(unsigned('0' & t(2 * INPUT_WIDTH downto INPUT_WIDTH + 1)) + unsigned('0' & b));	-- We should use an adder here
						t(INPUT_WIDTH - 1 downto 0) <= t(INPUT_WIDTH downto 1);
					else
						t(2 * INPUT_WIDTH downto 0) <= '0' & t(2 * INPUT_WIDTH downto 1);
					end if;
					ta <= '0' & ta(INPUT_WIDTH - 1 downto 1);

					if (counter = INPUT_WIDTH	) then
						counter <= counter;
					else
						counter <= counter + 1;
					end if;
				else -- We are in the done state
					ta <= ta;
					t <= t;
					counter <= counter;
				end if;
			end if;
		end process;
end architecture standard;